PK   ؐiV�n   ޾     cirkitFile.json�][����+�ΫZ�I��ɞ`a���HY,<�}����9�&N��_�u������	�̃=�,�ɯ?���ϓ���^������Ro���jr��t��o�O��*�N��n=�y�?L�>ǿ��o�uV�?>�W�j7o���+���3e��\�L������(��M��?Lo��q����UW��:T��K]{�\V7\eJy����,��f�*^��q���D˒嶬�2c܋L5�ʊRجvNȲ�L�+�8�e��2�0\9�p��L��g*uV��e��*ǥ��p]�8g��Fu9G>c\$L�M�YY�L2c��u�B��
�ȲlLc%�t�*j�9��橧U\��Hӑ)����gM �$������@NK	]�����&���0L>+rj�Ȝ�2����7J�I�4��aL��ej�Q�.��y�h�;���3��"/��
�p�#9�����d*�e]�,�_eʅi�M��Fs_��rf�іA=��]$��*q۶)\Q�<�uՄ9�)CmQdƸ�hH��l�����@��뵔�
l�]�8	�4��$r:U��T!�S��Nv���Nr:U���q�Bq�h:5/@��tj^�Nh��S���h:5-@��񦁓
��S^��̀>�x��9s�9�iܳ%�=`w��\�"��)J �M�T�0�3V)���`2�40P�h:�l #?���a�x��T��N�5*��Obn:�o�݈��8{���i�\/��6��o���	��B�E�h�$Z����W�Fhɣ��5�kZ�٨��B��A]ަa�U54��-|s++��~��m\�QC`��j��Q�� �54�F�"�!aA��BӨ�A�أ�V�Oā�[ָ=�����̺.6�K���u#F͞��9�D%��ž67@�(v�1�1j(6U�pC���8�N�n�Œ��+.V4\��<b.V4\�^�bh��2�����&4r|���A��t��^�����˼��^�rh��2�A���m��"/;�а��4DxyކF�.�4pwy��]^@A�i�Ws����  4�uy��X�ly� mw~Wc#H��i��Kd	�E�h�$Z�M�%'�bH�X-�uD�A/��/��/�0�A0��0��0�1�A��A� �`KKK"W�ŒŒŒŒŒŒŊŊŊŊ�#�A��A�z��^ˋ�� ᵼ8���E-�^ˋ�� ᵼh8����-�^ˋ��#Hx-/�� ᵼh8���rn˗i����>i��~��q;�|Zl���q�C_���zS՛��{��YL$�a��K�0��5�pM�v0M��X��s���_k�%f��i��k�YaL^3f�B�w�rPM'���ȏ��Qg,0`�i�;�������n�����llL.7��Auwb��o�@��c|�߃N��Q�C0+�������?�	��_Ucn��`�����_Ņl-x����O �T��d���"�ҧ�[�u�	,@z� m�Xo��&��M`�	�h����	� �_��kx��"�A�[���/�5�u�1@z� ��ߏ��><�XW>:�~S=-V�t������s�6�p��1����Y_!��}S��I��T�S�au��;;0�%\p�!
ll�=��Q��6��g�L���,�8�|�o�9�Ԧ��B�M3D)��X`9W�I˺K��6y� ��6a��h��b�����A�F�u���C��/K,��y�(_DB��!_�A�w��x�aOf���'@b�Ya�Ya�Ya�Y�=b,5+,5������H{��0���a��#����Ɇ0Jg��%(�~#Dp"�:pBbO&�=b]b1NQ��.e4W�w�Şu	��{�0����g�K0
8���.�w�ǁu_��g5�*F���meA����8�q�F�bFFPǧ8�'rM;��p����K��-^y�Q��
<���hu�"����5D����X�݇l�}�~`{��F�!��е�3�N��5�w�XC�*�P��*�P�+!�=��2�O�+�
��T��N��: �f��q�T� ��B�����z�:߿Ϲ�\�w(��T�� �Ƹ�ա��{�3.�u����j�Kpz���{�r^������4ء��z�/.3v�%���K�:J��� ���.�n������P;�6Q�e���}U�;�qi�C��nc�f.�v��^��K�� po��e�ׂ�פ��ϟݴ]<O��E���Z�1�B�_��Ml�W�E|X$EbX$ErX�EjX�EzX���a�9�a�=�a�;�A?�v?uǰ?��?��C��C��G��G��K��K�/a,�r9/6u���ob.s��/�]�X���>@��"SR���ȬԆ뢔N��<8���<��?9_��."6���li�����p�s{��f�Xov��]�~|\��"D����f��9���������|�����}��?�ϛwoߨ7�}��o���7�?���j���߶֟�_�Ghir�����z��b�(���ڦ���bS���.�R蟏~���r���7�L:;��o�z���ͻ�9�5X��b�~��}|Hg���S���Z���0����ַ��$�u�������W�9i���9�|!�mWߋ�v�W�(T0��7�0�~o���1\*�rYF�}�3��L��;�����T(](4V�Cᾌ��n{@nR�PpT�v����)�#��
�a���s�q�����p�#��
��E���Lb\��7��g�q�m���g�*���%�/���B��-ʤM��*L{��x��IU#��*sU9"9�R�۶IM��
�xAo���tW�I���bB��xU �u$<��4&9�Ҵ�-ҷu.1�BǮR%5<�+P���jRӈ�K�9�$�g�i�W唳��,7�8��VP���k}|��4	����qy�b]Bc�V��d��O|ƙ���u>S�q�����,v"�N�v�->���NP�����{�럎�z��.�	��<��W��<-voޮ��X'���y��N��uj��a��#~HS���Jd��U�%�ڶ��k�f���!�@=���F_�:��E|�UhU=_�g�:H��Cv*f���G��t)�g��Z!�<�@���4�V�R��:���l�M�Z/5�J��JS��+� V����~�!��gN*tjjf�_�_@��<�䀍�`� �9I,\@x ��~Q�0e��{���׏`�_�_3�O�az��~����x}\I��&�CJK���K�1�xƴr�e�s��A��������u���A	7 �U9�ς��:��	��v'�Q"ﰌF���qu��KO�d�����<w�(GŒ.��Bjq�O-�?a�Jހ0����NM�v>���%?MHǛ�4�K){�u�����WbaJ��`=����nF�K71J����:�w�&��O�%,f@Y\̴A々��ö]����C0�E�č��Ӫjѱ[�N�d\��b��lw��C�M����v�2 4?s�Ց)?ԋ�?DY#t\��WT���DL��出����nS�v����?�w|aP�G�|?i_;y?��?~��~2�(�ݻ��m�ݜ��*�W�EU��V����Ҷ��[B�׋���}h�}�������w������ƫw��g��6<�n���O��ʹ��R_Ί��P���q��h�urB�������K@ip��kQN�N����c��%�u���^θ.�`bّQ@:n�\)���p��t���p�p��2\W.��Hʻ���e\�Q�����倀�ːp�p�p�p�F� �u��ی:��8g��>�r�)5~��p�p�>�ܭ>�=����q�P�(A�23��i?^_%�R��7�������᮰�
p�&�k'�3��'�Z&��}�sF�urǜ}@��R�p������!�M������y��4�=!�`���(��K�1�t����U�d1g�S9�3c���͌�-H���q��"		7>�3�P�,L�0'(�����)�F��b�{���u�����p���8�\B0��lL h�������;'�Z8�º� �qo�����ɚ �����?W������Оs�w�Ξs)f�J���<P1��IHu.�X>�����(�\N�($>�|s���"\�~�mdW� ��Nz���xr-��Jb�t��*1 �JaK� !;�M�+�W�F���V�tYh|9Г2������PT,����g�/<m㠳1�|=a�L#�v6>�w%Ժ9b�|�O�K�o]vק �Q�'^'�3��JA�D�[�`vE�
ӨPv�F�)Qh��e	u���\�{�T.	�C�D^'�G����+��Zhybj4��u3&� i&\E	�}!F��}!vD$�@rf|��n�*�d�����Ā^Vne%��H���튘�����G7�:���&��DP>W��IX8(F�⁓;��2�G���S���,�q���k��{�!X,�)��n�0�����@��#3�����w~Wo~���E�n�?�WW��Փ_~���vW�ƞ|�2���PK
   ؐiV�n   ޾                   cirkitFile.jsonPK      =   8    